This is a resistive divider circuit.

R1 net_a net_b 10k
R2 net_b gnd 10k

*voltage supply
v1	net_a gnd sin (0 1V 10k) 	*sin (vdc vac_peak freq delay)  
	
.control
tran 2u 1ms
plot v(net_b) v(net_a)
.endc
.end
