Transient Analysis of Common source amplifier with Resistive load

.include spice_model.txt

M1 net_d net_g gnd gnd cmosn W=1u L=0.18u 
R1 net_d Vdd 10k

*voltage supply
V1 Vdd gnd dc 1.8
Vgs	net_g gnd sin (0.75 10mV 10k)	*sin (vdc vac_peak freq delay)

.control
tran 0.2u 1ms	
plot v(net_d) 
plot v(net_g)
.endc
.end
