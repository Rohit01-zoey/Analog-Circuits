DC Analysis of Common source amplifier with Resistive load

.include spice_model.txt

M1 net_d net_g gnd gnd cmosn W=1u L=0.18u 
R1 net_d Vdd 10k

*voltage supply
V1 Vdd gnd dc 1.8
Vgs	net_g gnd dc 0.75	

.control
save all @M1[vth]
save all @M1[gm]

dc Vgs 0 1.8 0.01
*plot v(net_d)  
*plot -i(V1)

*plot @M1[vth]
plot @M1[gm]
.endc
.end
