****************DEMO*****************
**********including the model file
.include cmos_130nm.txt
****************************
VDD net1 GND 1.5
RD net1 vout 10k
VG vin GND 0.6

* Mosfet M1  Drain Gate Source Body

M1 vout vin GND  GND NMOS W = 1u L = 130n
*******************ANALYSIS*************8
.control
*********DC Analysis
op
print @M1[id]

.endc
.end